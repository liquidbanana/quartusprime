LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LAB10PART4 IS
	PORT(CLOCK_50: IN STD_LOGIC;
	HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX2: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	HEX3: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END LAB10PART4;


ARCHITECTURE BEHAVIOR OF LAB10PART4 IS

	SIGNAL CLK: STD_LOGIC_VECTOR(0 TO 24);
	SIGNAL COUNT: STD_LOGIC_VECTOR(0 TO 1);
	
BEGIN

	PROCESS(CLOCK_50)
	BEGIN
	IF (CLOCK_50'EVENT AND CLOCK_50 = '1') THEN
		CLK <= CLK + 1;
		
		IF (CLOCK_50'EVENT AND CLOCK_50 = '1') THEN
			IF (CLK=0) THEN
				COUNT <= COUNT + 1;
			--ELSIF (COUNT = "11") THEN
				--COUNT <= "00";
				
			END IF;
		END IF;	
	END IF;
	END PROCESS;

	
	HEX3 <=	"0100001" WHEN COUNT = "00" ELSE
				"1000000" WHEN COUNT = "01" ELSE
				"1111001" WHEN COUNT = "10" ELSE
				"0000110"; --WHEN COUNT = "11";
				
				
	HEX2 <=	"0000110" WHEN COUNT = "00" ELSE
				"0100001" WHEN COUNT = "01" ELSE
				"1000000" WHEN COUNT = "10" ELSE
				"1111001"; --WHEN COUNT = "11";	
				
	
	HEX1 <=	"1111001" WHEN COUNT = "00" ELSE
				"0000110" WHEN COUNT = "01" ELSE
				"0100001" WHEN COUNT = "10" ELSE
				"1000000";-- WHEN COUNT = "11";
				
	HEX0 <=	"1000000" WHEN COUNT = "00" ELSE
				"1111001" WHEN COUNT = "01" ELSE
				"0000110" WHEN COUNT = "10" ELSE
				"0100001";-- WHEN COUNT = "11";			
					
				
END BEHAVIOR;