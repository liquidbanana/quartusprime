LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY part3 IS
PORT ( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
LEDR: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);
HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
HEX2: OUT STD_LOGIC_VECTOR(0 TO 6);
HEX3: OUT STD_LOGIC_VECTOR(0 TO 6);
HEX4: OUT STD_LOGIC_VECTOR(0 TO 6);
HEX5: OUT STD_LOGIC_VECTOR(0 TO 6));
END part3;

ARCHITECTURE struct OF part3 IS
	
	COMPONENT MUX
	PORT (S, U, V, W, X, Y, Z: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	M: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END COMPONENT;
	
	
	COMPONENT HEXDECODER
	PORT (C: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	D: OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	
	
	SIGNAL M0: STD_LOGIC_VECTOR(2 DOWNTO 0); 
	SIGNAL M1: STD_LOGIC_VECTOR(2 DOWNTO 0); 
	SIGNAL M2: STD_LOGIC_VECTOR(2 DOWNTO 0); 
	SIGNAL M3: STD_LOGIC_VECTOR(2 DOWNTO 0); 
	SIGNAL M4: STD_LOGIC_VECTOR(2 DOWNTO 0); 
	SIGNAL M5: STD_LOGIC_VECTOR(2 DOWNTO 0); 
	


BEGIN

	LEDR <= SW;
	
	U0: MUX PORT MAP(SW(9 DOWNTO 7), -- 000
	"000",
	"101",
	"100",
	"011",
	"010",
	"001",
	M0);
	
	
	
	U1: MUX PORT MAP(SW(9 DOWNTO 7), -- 001
	"001",
	"000",
	"101",
	"100",
	"011",
	"010",

	M1);
	

	U2: MUX PORT MAP(SW(9 DOWNTO 7),
	"010",
	"001",
	"000",
	"101",
	"100",
	"011",
	M2);
	

	U3: MUX PORT MAP(SW(9 DOWNTO 7),
	"011",
	"010",
	"001",
	"000",
	"101",
	"100",

	M3);
	

	U4: MUX PORT MAP(SW(9 DOWNTO 7),
	"100",
	"011",
	"010",
	"001",
	"000",
	"101",

	M4);
	
	
	U5: MUX PORT MAP(SW(9 DOWNTO 7),
	"101",
	"100",
	"011",
	"010",
	"001",
	"000",

	M5);

	
	H0: HEXDECODER PORT MAP(M0, HEX0);
	H1: HEXDECODER PORT MAP(M1, HEX1);
	H2: HEXDECODER PORT MAP(M2, HEX2);
	H3: HEXDECODER PORT MAP(M3, HEX3);
	H4: HEXDECODER PORT MAP(M4, HEX4);
	H5: HEXDECODER PORT MAP(M5, HEX5);
	
	
	
END struct;

