LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY MUX IS
PORT (S, U, V, W, X, Y, Z: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	M: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END MUX;


ARCHITECTURE MUX1 OF MUX IS

	SIGNAL NOT0_NOT1_NOT2: STD_LOGIC;
	SIGNAL NOT0_NOT1: STD_LOGIC;
	SIGNAL NOT0_NOT2: STD_LOGIC;
	SIGNAL NOT1_NOT2: STD_LOGIC; 
	SIGNAL NOT1: STD_LOGIC;
	SIGNAL NOT2: STD_LOGIC;


BEGIN 
	
	NOT0_NOT1_NOT2 <= NOT(S(0)) AND NOT(S(1)) AND NOT (S(2));
	NOT0_NOT1 <= NOT(S(0)) AND NOT(S(1)) AND S(2);
	NOT0_NOT2 <= NOT(S(0)) AND NOT (S(2)) AND S(1);
	NOT1_NOT2 <= NOT(S(1)) AND NOT (S(2)) AND S(0);
	NOT1 <= NOT(S(1)) AND S(0) AND S(2);
	NOT2 <= NOT(S(2)) AND S(0) AND S(1);

	
	M(2) <= 
	((NOT0_NOT1_NOT2 AND U(2))
	OR (NOT1_NOT2 AND V(2))
	OR (NOT0_NOT2 AND W(2))
	OR (NOT2 AND X(2))
	OR (NOT0_NOT1 AND Y(2))
	OR (NOT1 AND Z(2)));


	M(1) <= 
	((NOT0_NOT1_NOT2 AND U(1))
	OR (NOT1_NOT2 AND V(1))
	OR (NOT0_NOT2 AND W(1))
	OR (NOT2 AND X(1))
	OR (NOT0_NOT1 AND Y(1))
	OR (NOT1 AND Z(1)));


	M(0) <= 
	((NOT0_NOT1_NOT2 AND U(0))
	OR (NOT1_NOT2 AND V(0))
	OR (NOT0_NOT2 AND W(0))
	OR (NOT2 AND X(0))
	OR (NOT0_NOT1 AND Y(0))
	OR (NOT1 AND Z(0)));

END MUX1;