LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY LAB8PART3 IS 
	PORT (CLK, D: IN STD_LOGIC;
			Q: OUT STD_LOGIC);
			
			-- SW0 D INPUT
			-- SW1 CLK INPUT
			-- LEDR Q OUTPUT

END LAB8PART3;


ARCHITECTURE BEHAVIOR OF LAB8PART3 IS

	SIGNAL S, R, CLK1, S_G, R_G, QM, QB, D1, S1, R1, S_G1, R_G1, QS, QB2: STD_LOGIC;
	ATTRIBUTE KEEP: BOOLEAN;
	ATTRIBUTE KEEP OF S_G, R_G, QM, QB, S_G1, R_G1, QS, QB2: SIGNAL IS TRUE;

BEGIN
	S <= D;
	R <= NOT(D);
	
	CLK1 <= NOT(CLK);

	R_G <= (R) NAND CLK1;
	S_G <= S NAND CLK1;
	
	QM <= S_G NAND QB;
	QB <= R_G NAND QM;
	
	D1 <= QM;
	S1 <= D1;
	R1 <= NOT(D1);
	
	S_G1 <= S1 NAND CLK;
	R_G1 <= R1 NAND CLK;
	
	QS <= S_G1 NAND QB2;
	QB2 <= R_G1 NAND QS;

	Q <= QS;
END BEHAVIOR;