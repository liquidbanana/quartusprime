LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY TFLIPFLOP IS
	PORT(T, CLOCK, CLEAR: IN STD_LOGIC;
			Q: OUT STD_LOGIC);
END TFLIPFLOP;

ARCHITECTURE BEHAVIOR OF TFLIPFLOP IS
	SIGNAL TEMP: STD_LOGIC := '0';
BEGIN

	PROCESS(CLOCK)
	BEGIN
	IF (CLOCK'EVENT AND CLOCK='1') THEN 
		IF (CLEAR = '0') THEN
			TEMP <= '0';
		ELSIF (T = '1') THEN
			TEMP <= NOT(TEMP);
		END IF;
	END IF;
	END PROCESS;
	
	Q <= TEMP;
	
END BEHAVIOR;
