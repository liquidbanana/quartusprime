LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY LAB10PART2 IS
	PORT(SW1, SW0, CLOCK: IN STD_LOGIC;
	HEX0, HEX1, HEX2, HEX3: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));

END LAB10PART2;
ARCHITECTURE BEHAVIOR OF LAB10PART2 IS

	COMPONENT DECODER
	PORT (W, X, Y, Z: IN STD_LOGIC;
	DISP: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));	
	END COMPONENT;

	SIGNAL FLIP: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
	

BEGIN
	
	PROCESS(CLOCK, SW1)
	BEGIN
	IF (CLOCK'EVENT AND CLOCK = '1') THEN
		IF (SW0 = '0') THEN
			FLIP <= (OTHERS => '0');
		ELSIF (SW1 = '1') THEN
			FLIP <= FLIP + 1;
		END IF;
	END IF;
	END PROCESS;

	D0:DECODER PORT MAP(W => FLIP(3), X => FLIP(2), Y=> FLIP(1), Z=> FLIP(0), DISP => HEX0);
	D1:DECODER PORT MAP(W => FLIP(7), X => FLIP(6), Y=> FLIP(5), Z=> FLIP(4), DISP => HEX1);
	D2:DECODER PORT MAP(W => FLIP(11), X => FLIP(10), Y=> FLIP(9), Z=> FLIP(8), DISP => HEX2);
	D3:DECODER PORT MAP(W => FLIP(15), X => FLIP(14), Y=> FLIP(13), Z=> FLIP(12), DISP => HEX3);

END BEHAVIOR;