LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY COMPARATOR IS
	
	

END COMPARATOR;


ARCHITECTURE BEHAVIOR OF COMPARATOR IS

	

BEGIN 





END BEHAVIOR;