LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY CIRCB IS
	PORT (R,S,T,U: IN STD_LOGIC;
	ROUT, SOUT, TOUT, UOUT: OUT STD_LOGIC);

END CIRCB;

ARCHITECTURE BEHAVIOR OF CIRCB IS

	
BEGIN 

	ROUT <= NOT(R) AND NOT(S) AND T;
	SOUT <= NOT(R) AND NOT(S) AND NOT(T);
	TOUT <= NOT(R) AND NOT(S) AND NOT(T);
	UOUT <= NOT(R) AND NOT(S) AND U;


END BEHAVIOR;