LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY CIRCA IS
	PORT (R,S,T,U: IN STD_LOGIC;
	ROUT, SOUT, TOUT, UOUT: OUT STD_LOGIC);

END CIRCA;

ARCHITECTURE BEHAVIOR OF CIRCA IS
BEGIN 

		ROUT <= '0';
		SOUT <= R AND S AND T;
		TOUT <= R AND S AND NOT(T);
		UOUT <= (R AND S AND U) OR (R AND T AND U);



END BEHAVIOR;