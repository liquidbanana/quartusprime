LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
ENTITY DECODER IS
	PORT (BITS: IN STD_LOGIC_VECTOR(0 TO 3);
	HEXDISPLAY: OUT STD_LOGIC_VECTOR(0 TO 6));
END DECODER;
ARCHITECTURE BEHAVIOR OF DECODER IS
BEGIN 
	PROCESS(BITS)
	BEGIN
	CASE BITS IS
		WHEN "0000" => HEXDISPLAY <= "1000000"; -- 0
		WHEN "0001" => HEXDISPLAY <= "1111001"; -- 1
		WHEN "0010" => HEXDISPLAY <= "0100100"; -- 2
		WHEN "0011" => HEXDISPLAY <= "0110000"; -- 3		
		WHEN "0100" => HEXDISPLAY <= "0011001"; -- 4
		WHEN "0101" => HEXDISPLAY <= "0010010"; -- 5
		WHEN "0110" => HEXDISPLAY <= "0000010"; -- 6
		WHEN "0111" => HEXDISPLAY <= "1111000"; -- 7
		WHEN "1000" => HEXDISPLAY <= "0000000"; -- 8
		WHEN "1001" => HEXDISPLAY <= "0010000"; -- 9
		WHEN "1010" => HEXDISPLAY <= "0001000"; -- A
		WHEN "1011" => HEXDISPLAY <= "0000011"; -- B
		WHEN "1100" => HEXDISPLAY <= "1000110"; -- C
		WHEN "1101" => HEXDISPLAY <= "0100001"; -- D
		WHEN "1110" => HEXDISPLAY <= "0000110"; -- E
		WHEN "1111" => HEXDISPLAY <= "0001110"; -- F
		WHEN OTHERS => HEXDISPLAY <= "1111111"; -- OTHER
	END CASE;
	END PROCESS;
END BEHAVIOR;