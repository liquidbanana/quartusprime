LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LAB10PART3 IS
	PORT(CLOCK_50: IN STD_LOGIC;
	HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END LAB10PART3;


ARCHITECTURE BEHAVIOR OF LAB10PART3 IS

	COMPONENT DECODER IS
	PORT (BITS: IN STD_LOGIC_VECTOR(0 TO 3);
	HEXDISPLAY: OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	
	SIGNAL CLK: STD_LOGIC_VECTOR(0 TO 24);
	SIGNAL COUNT: STD_LOGIC_VECTOR(0 TO 3);
	
	
BEGIN

	PROCESS(CLOCK_50)
	BEGIN
	IF (CLOCK_50'EVENT AND CLOCK_50 = '1') THEN
		CLK <= CLK + 1;
		IF (CLOCK_50'EVENT AND CLOCK_50 = '1') THEN
			IF (CLK=0) THEN
				COUNT <= COUNT + 1;
			ELSIF (COUNT = "1010") THEN
				COUNT <= "0000";
			END IF;
		END IF;	
	END IF;
	END PROCESS;
	h0: DECODER PORT MAP(BITS => COUNT, HEXDISPLAY => HEX0);
	
END BEHAVIOR;