LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY HEXADECIMALDECODER IS

		PORT (W, X, Y, Z: IN STD_LOGIC;
				HEXDISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
				
END HEXADECIMALDECODER;

ARCHITECTURE DECODER OF HEXADECIMALDECODER IS
	
BEGIN 
	
	HEXDISPLAY(0) <= (NOT(W) AND NOT(X) AND NOT(Y) AND Z) OR (NOT(W) AND X AND NOT(Y) AND NOT(Z)) OR (W AND X AND NOT(Y) AND Z) OR (W AND NOT(X) AND Y AND Z);
	HEXDISPLAY(1) <= (NOT(W) AND X AND NOT(Y) AND Z) OR (W AND X AND NOT(Z)) OR (W AND Y AND Z)  OR (X AND Y AND  NOT(Z));
	HEXDISPLAY(2) <= (NOT(W) AND NOT(X) AND Y AND NOT(Z)) OR (W AND X AND NOT(Z)) OR (W AND X AND Y);
	HEXDISPLAY(3) <= (NOT(W) AND NOT(X) AND NOT(Y) AND Z) OR (NOT(W) AND X AND NOT(Y) AND NOT(Z)) OR (X AND Y AND Z) OR (W AND NOT(X) AND Y AND NOT(Z));
	HEXDISPLAY(4) <= (NOT(W) AND Z) OR (NOT(W) AND X AND NOT(Y)) OR (NOT(X) AND NOT(Y) AND Z);
	HEXDISPLAY(5) <= (NOT(W) AND NOT(X) AND Z) OR (NOT(W) AND NOT(X) AND Y) OR (NOT(W) AND Y AND Z) OR (W AND X AND NOT(Y) AND Z); 
	HEXDISPLAY(6) <= (NOT(W) AND NOT(X) AND NOT(Y)) OR (W AND X AND NOT(Y) AND NOT(Z)) OR (NOT(W) AND X AND Y AND Z);

END DECODER;
