LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY LAB10PART11 IS

	PORT(SW1, SW0, CLK: IN STD_LOGIC;
			QOUTBAR: OUT STD_LOGIC;
			HEX0, HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO  0));

END LAB10PART11;

ARCHITECTURE BEHAVIOR OF LAB10PART11 IS

	COMPONENT TFLIPFLOP
	PORT(T, CLOCK, CLEAR: IN STD_LOGIC;
			Q: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT HEXADECIMALDECODER
	PORT (W, X, Y, Z: IN STD_LOGIC;
			HEXDISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));		
	END COMPONENT;
	
	SIGNAL ENABLE: STD_LOGIC;
	SIGNAL CLR: STD_LOGIC;
	
	SIGNAL Q0: STD_LOGIC;
	SIGNAL Q1: STD_LOGIC;
	SIGNAL Q2: STD_LOGIC;
	SIGNAL Q3: STD_LOGIC;
	SIGNAL Q4: STD_LOGIC;
	SIGNAL Q5: STD_LOGIC;
	SIGNAL Q6: STD_LOGIC;
	SIGNAL Q7: STD_LOGIC;
	
	SIGNAL Q1IN: STD_LOGIC;
	SIGNAL Q2IN: STD_LOGIC;
	SIGNAL Q3IN: STD_LOGIC;
	SIGNAL Q4IN: STD_LOGIC;
	SIGNAL Q5IN: STD_LOGIC;
	SIGNAL Q6IN: STD_LOGIC;
	SIGNAL Q7IN: STD_LOGIC;
	
BEGIN
	
	Q1IN <= Q0 AND SW1;
	Q2IN <= Q1IN AND Q1;
	Q3IN <= Q2IN AND Q2;
	Q4IN <= Q3IN AND Q3;
	Q5IN <= Q4IN AND Q4;
	Q6IN <= Q5IN AND Q5;
	Q7IN <= Q6IN AND Q6;
	
	Q0CALL: TFLIPFLOP PORT MAP(T => SW1, CLOCK => CLK, CLEAR => SW0, Q => Q0);
	Q1CALL: TFLIPFLOP PORT MAP(T => Q1IN, CLOCK => CLK, CLEAR => SW0, Q => Q1);
	Q2CALL: TFLIPFLOP PORT MAP(T => Q2IN, CLOCK => CLK, CLEAR => SW0, Q => Q2);
	Q3CALL: TFLIPFLOP PORT MAP(T => Q3IN, CLOCK => CLK, CLEAR => SW0, Q => Q3);
	Q4CALL: TFLIPFLOP PORT MAP(T => Q4IN, CLOCK => CLK, CLEAR => SW0, Q => Q4);
	Q5CALL: TFLIPFLOP PORT MAP(T => Q5IN, CLOCK => CLK, CLEAR => SW0, Q => Q5);
	Q6CALL: TFLIPFLOP PORT MAP(T => Q6IN, CLOCK => CLK, CLEAR => SW0, Q => Q6);
	Q7CALL: TFLIPFLOP PORT MAP(T => Q7IN, CLOCK => CLK, CLEAR => SW0, Q => Q7);
	
	H0: HEXADECIMALDECODER PORT MAP(W => Q3, X => Q2, Y => Q1, Z => Q0, HEXDISPLAY => HEX0);
	H1: HEXADECIMALDECODER PORT MAP(W => Q7, X => Q6, Y => Q5, Z => Q4, HEXDISPLAY => HEX1);
	
END BEHAVIOR;




