LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY LAB74 IS
	PORT (SW: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
	LEDR: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
	HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
	--HEX2: OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX3: OUT STD_LOGIC_VECTOR(0 TO 6);
	--HEX4: OUT STD_LOGIC_VECTOR(0 TO 6);
	HEX5: OUT STD_LOGIC_VECTOR(0 TO 6));
	
END LAB74;


ARCHITECTURE BEHAVIOR OF LAB74 IS

	COMPONENT DECODER IS
	PORT (A,B,C,D: IN STD_LOGIC;
	HEXDISPLAY: OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;

	COMPONENT FULLADDER IS
	PORT (A, B, C: IN STD_LOGIC;
		S, C0: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT MUX
	PORT (I0, I1, S: IN STD_LOGIC;
	MUXOUT: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT CIRCA
	PORT (R,S,T,U: IN STD_LOGIC;
	ROUT, SOUT, TOUT, UOUT: OUT STD_LOGIC);
	END COMPONENT;

	COMPONENT CIRCB
	PORT (R,S,T,U: IN STD_LOGIC;
	ROUT, SOUT, TOUT, UOUT: OUT STD_LOGIC);
	END COMPONENT;
	

	SIGNAL S3: STD_LOGIC;
	SIGNAL S2: STD_LOGIC;
	SIGNAL S1: STD_LOGIC;
	SIGNAL S0: STD_LOGIC;
	
	SIGNAL C1: STD_LOGIC;
	SIGNAL C2: STD_LOGIC;
	SIGNAL C3: STD_LOGIC;
	SIGNAL Cout: STD_LOGIC;
	
	
	SIGNAL COMP3: STD_LOGIC;
	SIGNAL COMP2: STD_LOGIC;
	SIGNAL COMP1: STD_LOGIC;
	SIGNAL COMP0: STD_LOGIC;
	SIGNAL COMPARATOR: STD_LOGIC;
	
	SIGNAL A3OUT: STD_LOGIC;
	SIGNAL A2OUT: STD_LOGIC;
	SIGNAL A1OUT: STD_LOGIC;
	SIGNAL A0OUT: STD_LOGIC;
	
	SIGNAL B3OUT: STD_LOGIC;
	SIGNAL B2OUT: STD_LOGIC;
	SIGNAL B1OUT: STD_LOGIC;
	SIGNAL B0OUT: STD_LOGIC;
	
	SIGNAL COMP7: STD_LOGIC;
	SIGNAL COMP6: STD_LOGIC;
	SIGNAL COMP5: STD_LOGIC;
	SIGNAL COMP4: STD_LOGIC;
	
	SIGNAL COMP11: STD_LOGIC;
	SIGNAL COMP10: STD_LOGIC;
	SIGNAL COMP9: STD_LOGIC;
	SIGNAL COMP8: STD_LOGIC;
	

BEGIN 
	
	-- HEX 5, 3
	H5: DECODER PORT MAP(A => SW(7), B => SW(6), C => SW(5), D => SW(4), HEXDISPLAY => HEX5);
	H3: DECODER PORT MAP(A => SW(3), B => SW(2), C => SW(1), D => SW(0), HEXDISPLAY => HEX3);
	
	-- HEX 1
	F0: FULLADDER PORT MAP(A => SW(4), B => SW(0), C => SW(8), S => S0, C0 => C1);
	F1: FULLADDER PORT MAP(A => SW(5), B => SW(1), C => C1, S => S1, C0 => C2);
	F2: FULLADDER PORT MAP(A => SW(6), B => SW(2), C => C2, S => S2, C0 => C3);
	F3: FULLADDER PORT MAP(A => SW(7), B => SW(3), C => C3, S => S3, C0 => Cout);
	
	
	M3: MUX PORT MAP(I0 => S3, I1 => '1', S => Cout, MUXOUT => COMP3);
	M2: MUX PORT MAP(I0 => S2, I1 => '1', S => Cout, MUXOUT => COMP2);
	M1: MUX PORT MAP(I0 => S1, I1 => '1', S => Cout, MUXOUT => COMP1);
	M0: MUX PORT MAP(I0 => S0, I1 => '1', S => Cout, MUXOUT => COMP0);

	COMPARATOR <= (COMP3 AND COMP2) OR (COMP3 AND COMP1);
	HEX1(0) <= COMPARATOR;
	HEX1(1) <= '0';
	HEX1(2) <= '0';
	HEX1(3) <= COMPARATOR;
	HEX1(4) <= COMPARATOR;
	HEX1(5) <= COMPARATOR;
	HEX1(6) <= '1';

	
	-- HEX 1
	A0: CIRCA PORT MAP(R => S3, S => S2, T => S1, U => S0, ROUT => A3OUT, SOUT => A2OUT, TOUT => A1OUT, UOUT => A0OUT);
	B0: CIRCB PORT MAP(R => S3, S => S2, T => S1, U => S0, ROUT => B3OUT, SOUT => B2OUT, TOUT => B1OUT, UOUT => B0OUT);
	
	M7: MUX PORT MAP(I0 => A3OUT, I1 => B3OUT, S => Cout, MUXOUT => COMP7);
	M6: MUX PORT MAP(I0 => A2OUT, I1 => B2OUT, S => Cout, MUXOUT => COMP6);
	M5: MUX PORT MAP(I0 => A1OUT, I1 => B1OUT, S => Cout, MUXOUT => COMP5);
	M4: MUX PORT MAP(I0 => A0OUT, I1 => B0OUT, S => Cout, MUXOUT => COMP4);
	
	
	M11: MUX PORT MAP(I0 => S3, I1 => COMP7, S => COMPARATOR, MUXOUT => COMP11);
	M10: MUX PORT MAP(I0 => S2, I1 => COMP6, S => COMPARATOR, MUXOUT => COMP10);
	M9: MUX PORT MAP(I0 => S1, I1 => COMP5, S => COMPARATOR, MUXOUT => COMP9);
	M8: MUX PORT MAP(I0 => S0, I1 => COMP4, S => COMPARATOR, MUXOUT => COMP8);
	
	
	H1: DECODER PORT MAP(A => COMP11, B => COMP10, C => COMP9, D => COMP8, HEXDISPLAY => HEX0);


END BEHAVIOR;







	
	
	
	

