LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY lab7part2 IS 
PORT (SW: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		LEDR: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX1: OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX2: OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX3: OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX4: OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX5: OUT STD_LOGIC_VECTOR(0 TO 6));	

END lab7part2;

ARCHITECTURE behavior OF lab7part2 IS
		SIGNAL A3: STD_LOGIC;
		SIGNAL A2: STD_LOGIC;
		SIGNAL A1: STD_LOGIC;
		SIGNAL A0: STD_LOGIC;
		SIGNAL Z: STD_LOGIC;
		SIGNAL M3: STD_LOGIC;
		SIGNAL M2: STD_LOGIC;
		SIGNAL M1: STD_LOGIC;
		SIGNAL M0: STD_LOGIC;
		

BEGIN
		
	--	A3 <= NOT((NOT(SW(3)) AND NOT(SW(2))) OR (NOT(SW(3)) AND SW(1)));
		A3 <= '0';
		A2 <= SW(3) AND SW(2) AND SW(1);
		A1 <= SW(3) AND SW(2) AND NOT(SW(1));
		A0 <= (SW(3) AND SW(2) AND SW(0)) OR (SW(3) AND SW(1) AND SW(0));
		Z <= (SW(3) AND SW(2)) OR (SW(3) AND SW(1));
		
	
		M3 <= (NOT(Z) AND SW(3)) OR (A3 AND Z);
		M2 <= (NOT(Z) AND SW(2)) OR (A2 AND Z);
		M1 <= (NOT(Z) AND SW(1)) OR (A1 AND Z);
		M0 <= (NOT(Z) AND SW(0)) OR (A0 AND Z);
		
		HEX1(0) <= Z;
		HEX1(1) <= '0';
		HEX1(2) <= '0';
		HEX1(3) <= Z;
		HEX1(4) <= Z;
		HEX1(5) <= Z;
		HEX1(6) <= '1';
		
		
		HEX0(0) <= (NOT(M3) AND M2 AND NOT(M1) AND NOT(M0)) OR (NOT(M3) AND NOT(M2) AND NOT(M1) AND M0);
		HEX0(1) <= (NOT(M3) AND M2 AND NOT(M1) AND M0) OR (NOT(M3) AND M2 AND M1 AND NOT(M0));
		HEX0(2) <= (NOT(M3) AND NOT(M2) AND M1 AND NOT(M0));
		HEX0(3) <= (NOT(M3) AND NOT(M2) AND NOT(M1) AND M0) OR (NOT(M3) AND M2 AND NOT(M1) 
		AND NOT(M0)) OR (NOT(M3) AND M2 AND M1 AND M0);
		HEX0(4) <= (NOT(M3) AND M0) OR (NOT(M3) AND M2 AND NOT(M1)) OR (NOT(M2) AND NOT(M1) AND M0);
		HEX0(5) <= (NOT(M3) AND NOT(M2) AND M0) OR (NOT(M3) AND NOT(M2) AND M1) OR (NOT(M3) AND M1 AND M0);
		HEX0(6) <= (NOT(M3) AND NOT(M2) AND NOT(M1)) OR (NOT(M3) AND M2 AND M1 AND M0);
		
	

END behavior;
