LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY LAB10PART1 IS
	PORT(CLK: IN STD_LOGIC;
			SW: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			QOUTBAR: OUT STD_LOGIC;
			HEX0, HEX1: OUT STD_LOGIC_VECTOR(6 DOWNTO  0));

END LAB10PART1;
------------------------------------------------------------------------------------------------------

ARCHITECTURE BEHAVIOR OF LAB10PART11 IS

	COMPONENT TFLIPFLOP
	PORT(T, CLOCK, CLEAR: IN STD_LOGIC;
			Q: OUT STD_LOGIC);
	END COMPONENT;
	
	COMPONENT DECODER
	PORT (W, X, Y, Z: IN STD_LOGIC;
			DISP: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));		
	END COMPONENT;
		
	SIGNAL Q0: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TEMP: STD_LOGIC_VECTOR(6 DOWNTO 0);
------------------------------------------------------------------------------------------------------
	
BEGIN
	
	TEMP(0) <= Q0(0) AND SW(1);
	TEMP(1) <= TEMP(0) AND Q0(1);
	TEMP(2) <= TEMP(1) AND Q0(2);
	TEMP(3) <= TEMP(2) AND Q0(3);
	TEMP(4) <= TEMP(3) AND Q0(4);
	TEMP(5) <= TEMP(4) AND Q0(5);
	TEMP(6) <= TEMP(5) AND Q0(6);
	
	TFF0: TFLIPFLOP PORT MAP(T => SW(1), CLOCK => CLK, CLEAR => SW(0), Q => Q0(0));
	TFF1: TFLIPFLOP PORT MAP(T => TEMP(0), CLOCK => CLK, CLEAR => SW(0), Q => Q0(1));
	TFF2: TFLIPFLOP PORT MAP(T => TEMP(1), CLOCK => CLK, CLEAR => SW(0), Q => Q0(2));
	TFF3: TFLIPFLOP PORT MAP(T => TEMP(2), CLOCK => CLK, CLEAR => SW(0), Q => Q0(3));
	TFF4: TFLIPFLOP PORT MAP(T => TEMP(3), CLOCK => CLK, CLEAR => SW(0), Q => Q0(4));
	TFF5: TFLIPFLOP PORT MAP(T => TEMP(4), CLOCK => CLK, CLEAR => SW(0), Q => Q0(5));
	TFF6: TFLIPFLOP PORT MAP(T => TEMP(5), CLOCK => CLK, CLEAR => SW(0), Q => Q0(6));
	TFF7: TFLIPFLOP PORT MAP(T => TEMP(6), CLOCK => CLK, CLEAR => SW(0), Q => Q0(7));
	
	H0: DECODER PORT MAP(W => Q0(3), X => Q0(2), Y => Q0(1), Z => Q0(0), DISP => HEX0);
	H1: DECODER PORT MAP(W => Q0(7), X => Q0(6), Y => Q0(5), Z => Q0(4), DISP => HEX1);
	
END BEHAVIOR;