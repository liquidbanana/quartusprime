LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;


ENTITY MUX IS
	PORT (I0, I1, S: IN STD_LOGIC;
	MUXOUT: OUT STD_LOGIC);
END MUX;


ARCHITECTURE BEHAVIOR OF MUX IS
BEGIN 
	MUXOUT <= (I0 AND NOT(S)) OR (I1 AND S);

END BEHAVIOR;