LIBRARY IEEE;
USE STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LAB7PART6 IS
	PORT (SW: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
			LEDR: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			HEX0: OUT STD_LOGIC_VECTOR(0 TO 6);
			HEX1: OUT STD_LOGIC_VECTOR(0 TO 6));

END LAB7PART6;

ARCHITECTURE BEHAVIOR OF LAB7PART6 IS

	COMPONENT DECODER
	PORT (HEXDIS1, HEXDIS0: IN STD_LOGIC;
	HEXDISPLAY: OUT STD_LOGIC_VECTOR(0 TO 6));
	END COMPONENT;
	
	SIGNAL HEXDIS0: STD_LOGIC_VECTOR(0 TO 6);
	SIGNAL HEXDIS1: STD_LOGIC_VECTOR(0 TO 6);s
	
	SIGNAL SWITCH_INPUT: INTEGER;
	SIGNAL TENSPLACE: INTEGER;
	SIGNAL ONESPLACE: INTEGER;

BEGINS
	SWITCH_INPUT <= to_integer(unsigned(SW(0 TO 5));
	PROCESS: PROCESS(SWITCH_INNPUT);
	IF SWITCH_INPUT > 59 THEN TENSPLACE <= 6;
	ONESPLACE <= SWITCH_INPUT - 60;
	ELSIF SWITCH_INPUT > 49 THEN TENSPLACE <= 5;
	ONESPLACE <= SWITCH_INPUT - 50;
	ELSIF SWITCH_INPUT > 39 THEN TENSPLACE <= 4;
	ONESPLACE <= SWITCH_INPUT - 40;
	ELSIF SWITCH_INPUT > 29 THEN TENSPLACE <=3;
	ONESPLACE <= SWITCH_INPUT - 30;
	ELSIF SWITCH_INPUT > 19 THEN TENSPLACE <= 2;
	ONESPLACE <= SWITCH_INPUT - 20;
	ELSIF SWITCH_INPUT > 9 THEN TENSPLACE <= 1;
	ONESPLACE <= SWITCH_INPUT - 10;
	ELSE TENSPLACE <= 0;
	END IF;
	END PROCESS;
	
	HEXDIS1 <= to_integer(unsigned(tensplace,6));
	HEXDIS0 <= to_integer(unsigned(onesplace,6));
	
	H1: DECODER PORT MAP(HEXDIS1, HEXDISPLAY => HEX1);
	H0: DECODER PORT MAP(HEXDIS0, HEXDISPLAY => HEX0);
	
	
END BEHAVIOR;